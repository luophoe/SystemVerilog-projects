///////////////////////////////////////////////////////////////////////////
// (c) Copyright 2013 Cadence Design Systems, Inc. All Rights Reserved.
//
// File name   : control.sv
// Title       : Control Module
// Project     : SystemVerilog Training
// Created     : 2013-4-8
// Description : Defines the Control module
// Notes       :
// 
///////////////////////////////////////////////////////////////////////////

// import SystemVerilog package for opcode_t and state_t

module control import typedefs::*; (
                output logic      load_ac ,
                output logic      mem_rd  ,
                output logic      mem_wr  ,
                output logic      inc_pc  ,
                output logic      load_pc ,
                output logic      load_ir ,
                output logic      halt    ,
                input  opcode_t opcode  , // opcode type name must be opcode_t
                input             zero    ,
                input             clk     ,
                input             rst_   
                );
// SystemVerilog: time units and time precision specification
timeunit 1ns;
timeprecision 100ps;
logic a, h, k, j, s;
state_t st;

always_ff @(posedge clk or negedge rst_)
  if (!rst_)
     st = st.first();    
  else
     st = st.next();
  
always_comb
  begin
   a = (opcode == 2 || opcode == 3 || opcode == 4 || opcode == 5) ? 1 : 0;
   h = (opcode == 0) ? 1 : 0;
   k = (opcode == 1 && zero) ? 1 : 0;
   j = (opcode == 7) ? 1 : 0;
   s = (opcode == 6) ? 1 : 0;

   unique case (st)
      3'b000   : begin mem_rd =  0; load_ir = 0; halt = 0; inc_pc = 0;load_ac = 0; load_pc = 0; mem_wr = 0; end
      3'b001   : begin mem_rd =  1; load_ir = 0; halt = 0; inc_pc = 0;load_ac = 0; load_pc = 0; mem_wr = 0; end
      3'b010   : begin mem_rd =  1; load_ir = 1; halt = 0; inc_pc = 0;load_ac = 0; load_pc = 0; mem_wr = 0; end
      3'b011   : begin mem_rd =  1; load_ir = 1; halt = 0; inc_pc = 0;load_ac = 0; load_pc = 0; mem_wr = 0; end
      3'b100   : begin mem_rd =  0; load_ir = 0; halt = h; inc_pc = 1;load_ac = 0; load_pc = 0; mem_wr = 0; end
      3'b101   : begin mem_rd =  a; load_ir = 0; halt = 0; inc_pc = 0;load_ac = 0; load_pc = 0; mem_wr = 0; end
      3'b110   : begin mem_rd =  a; load_ir = 0; halt = 0; inc_pc = k;load_ac = a; load_pc = j; mem_wr = 0; end
      3'b111   : begin mem_rd =  a; load_ir = 0; halt = 0; inc_pc = j;load_ac = a; load_pc = j; mem_wr = s; end
      default  : begin mem_rd =  0; load_ir = 0; halt = 0; inc_pc = 0;load_ac = 0; load_pc = 0; mem_wr = 0; end
   endcase
 end
 
endmodule
